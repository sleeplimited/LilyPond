BZh91AY&SYfz�B �߀Pyc����������P>)@��TRH�����S~��OT�RhyOI�D�d�m!�M21M0�&�F	���#C@p�L�FL0	��bd4���4�#��i�`��244D�e4�S��	
z����bf�M{9U�SB!�G�{�PZ� �Ʉ������|���MmUy�Z`�F!U���hcIV Vaנ_n�60�|�J#���&�1������.N�����q=$j�Hb�K�Ǜ����ccY��*k;��9a�x��97 )�,���'1��0��P8_��C6ړ&fM\x���x|_�y�4�
�h�h|�L{�	H7����NZ�]�.��j�u�IX<XH�SF{�d��f��v�s~z�i4J4f���/@�clc}Ͷ�m�pB�W?w2'�Lk��.lJ*Z�U�`��N��E�`:���eK�r��,���������֦��jc1�4�`��eL�3iQ�F/�|�ǆI�'u�n������)l��ӯ������������@��;`��-F�o�~w���k���T���/�Y>J6��ې�\�}�Wa�x�9�Ǽ;�~�"jYnZ�Bg]�����1���Ӗģ���K�����~/�f޷Ƅ{����0e퍦���K�#|�T�(!��alI���d�����u\��Bs�ڹ���e�T��R����Q��Q����9 ���s��B�S�����G2�LbRoy-X&*C�hʨt&a]�K�YU(.�����p�`o�J=�")�V�0}3�P&]�:6+"�KR;�z~��$�ͷ��eȆ�A��� ���7�9��*(��;��?�ZP�us�#-���[M�z����'�B%�.lq���U��-��	�[�p,���}%QƁ�7 (�F�&��$��2F
���i�	�tL���AP��ui(%T�A��,9;�'a=�I@PtQ`2*�$1�&��؜�͎�90��\� {��l5���B�0KB[B[e	��|�`��׀˩�,MC4��o��\��m}'A�ʔYl�Kʆ ��pyA�s��=�Ǯ�M�ϯl��)eˢKJ���-��E&y�"���oVa��2�QÎH,e%Jb��'���|^�]�*��S,�^<ID+Y���E
6�p�p�LE�+ *xqz���O��-��z�:�%��sd�l��Ă���`�%�FLM~�O�c
����"��.�p� ����